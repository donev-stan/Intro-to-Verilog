module my_or_gate (
  input A, B,
  output C
);
  
  assign C = A | B;
  
endmodule