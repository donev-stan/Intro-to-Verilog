module tb ();
  parameter N = 3;
  
  reg [(1<<N)-1:0] X;
  wire [N-1:0] Y;
  
  encoder 
  #(.N(N))
  u_encoder (
    .X(X),
    .Y(Y)
  );
  
  initial begin
    repeat (10)
      #10 X = $random();
    #10 $finish();
  end
  
  initial begin
    $dumpfile("dump.vcd"); $dumpvars;
  end
  
endmodule