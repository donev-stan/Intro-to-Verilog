module my_not_gate (
  input A,
  output C
);
  
  assign C = ~A;
  
endmodule