module my_xor_gate (
  input A, B,
  output C
);
  
  assign C = A ^ B;
  
endmodule